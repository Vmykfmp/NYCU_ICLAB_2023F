/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2023 Autumn IC Design Laboratory 
Lab09: SystemVerilog Design and Verification 
File Name   : PATTERN.sv
Module Name : PATTERN
Release version : v1.0 (Release Date: Nov-2023)
Author : Jui-Huang Tsai (erictsai.10@nycu.edu.tw)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/
`define PAT_NUM 100000
`include "Usertype_BEV.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
b\M^3.W^\XCcPS;+eVb06.I:bMB1A[<M5[RPI#IWIGbLKFF17U#b1)7RgVdL)_+-
N)+F_]<UH/\4<(5a[_CK808L)9e]@Z<SR6SM9&__+\./W5V[U[_7a1-;>:2J+f>I
cJ_DLg[7N2=5?R(8e:,[+)RP8K0c3XG0/]b701T>#.LgC\5[d)V\]a=ZbXPZ2.4Y
<WP+7d4NK[K>f(b>8>e^W:;QZ--@^^T8b7,c&eQe#&GZ8_#6KDRVBAQJ[OCX7\_M
13e)0#W@O@H2+OMbH>S#:E;?2DF\[#@d(dU:,?XZ0=bV2Y.];f5BgC9_??II?O3:
G0W>fUPW,F0gd,]7G<;?)0TI6bdCIGA5S;OXA6X_8HCDBHd1=.]YGM[T6Q-?W;Y:
R?08PXEOR_/XV59+M\f<X9L0.c]I</=&VVMUWF4;4-JRN^JH87MaT3XLN0@<)a7_
1AMP1c,>9+W-4@Q4AKaDX<c]:37SW6L/Z/X/1#Y<V4?SKZ52S1FfIP<gg[eGC.DX
02:>X=&eL>/=DD,STXN:-Y1g3F&V;MA,6ABaHA;>L#=L3f+8J\7]N\MDM&^6JCHC
3J2P)(+Ob0f,4R&\^3;7[OI0[g)g\3ER^S5?FD@ZHI[6N#?J;W^B:OE-a[A3UWYR
/7IU1a\UJ.[NWVD@@7<LI?EI;&]eQA^4c,a:08Y@?>F+G;^M8/d:-U3bc]@d>DO2
]0#L,(YG]SC-f:&a-bcAdZV0)W@NFaCD\BHcOW&_a.YGG+2>36NZgb;99DM&_[NR
KdME].1eCDPa;UQQAP:#_@IRKG&fFbQE^T_c^EMf7b?f6S>X,G78_gS8fO_FSUVX
S:DL>YW4H1<D](X?.F;)@Pc^b9<?BIZ7Zc?SN<PS47H+CMH,/-A>>E5.-0<K^YXE
c+&CK+[HdQ5Zd:YY4[=X9(]^N8,-Y0C@52SE@WI4S<d?@J][>V9(aD=F4I1JMUV7
]fb@G3#?)FGD.+OZ0ZIg\F3=Q_1D3\X9YQ2E0),U0M[Fc4O.1c]DN_\R&-D8=ES7
1@@3VRY(B>PTSIa>L/I/Q]<>/,c>CD6S.N_CdeLBcg_f4]I-b\HDO:a8D5XHOU@<
9.AC[M_R-ZT5]VB.\^[cR0T\42,-@4/)FJ:\+^A-D5&/R>][#]bAL?fOZ94=WP8Z
CUQ,P?K;1/+@S[)95]HfS\H(cg3Z7@Ua(R2WSaE(@<U=]Db[c,NY5cQS9?gYdE/W
Q)[-JdC[<g)[e8(,7XEGaIBLPB[(gHMd7N#9&(Z@;:28AU9,@9.HcVfJd>KHc#A,
8:^=<F5(WJ-QR\\]KMI2,C4?.OQGG0YQ@YVJ_c#OKF7YA6C<^c;[;#gO0VcAIadb
fGH1bd<F??.b?0Mc#\@9b+9/1AD9R<QfBJ.Z[UT2c1+7YHaN9O09TJ[YTR?RZY,-
d7IUJd?+LRYF#gcG?S[b3ZKT;0>Zg@8eZSP<S__CCEB-@BX)_.=/NE=^WW8f:ZXZ
[T-UV].35)dP.0e^Ja-(a-aG+1&P3P\>e218eCG/?<1Xb_/c2f9&447XE]0,fbdb
cRLg)(P#3DgG7=N?Ib4GX=[R;L([;2.+;P-W/&b/+0Mb6dL2c/37OTMcDa2&XYV9
X].8I4+4VeB:I]PE#IMYbZL&Y\R(P&FS8ETJ:1YLgH66WRNd[>Hd,4_aY6Y>_Zg?
U7<_(,Q^f_192N(0K(^]\Qg1&4JX)g&UVHKU9AI6(DTALLI^Y&=]Z+B_L4P8UHK)
)9L3Y9)d89Q>\dgD+^f3@U/2ebU\<.V^ZUXW6]c?FDdUZg=,:61-=V,9cD8>>M;N
0</7DSN5T@;GMIW^WZ]Z&<?G#be9;7^Yf88NZ/B8+S870R=5g<ELB(8EdG.38&7,
^MMXL8Bc7Ma0Y620I<A<BdVB.Z>NbJSSA,6:XO9L2Sg[^U:7]KLg/eDXRAML7g,_
3BZ(2;:UKfed,+BcfXN#K;Z9FC1B59I)=aJ9UB^e1g8FD^,<NJ0<M(KZ\f)65E12
[V0HA(c8g<6,=b^8CMO7PW1_\e4G^\A63-SV):+[>R/8TMZEd.L?+VeH]9H6_E\&
W2=72Nf_L#PZ4NZ+;UVe363_&OY3LdABW0eGK/7-W-3eJX]cSAZ;AO-b(X+a,f1>
>&//GRY>DP3d7Z^,#ME>.<&#2T8M:Y30-1=LW2G9&\b+80]BH&,GL7a.?.3ZI_gC
@6d>8-Y5?+]S+??U0M9eZ0L#IF+<f/3)aFc8T\(+g>G]@#8:G;DO5O)gaG.ZUD@R
CN-+)V:NOGBC:#3L]TJWDC,BPE32X-1K1f-4)eAJRK6/GY(^UWSa^>.>_2>,1D@H
/+&S@U:1GCVXJdQae8?gZg_XKeJRM&Wg&X#[]QGf-]CH&<_3[9I.fV_.?F24,DWA
afVNX26^(8fWZFI8].&NX_?1A.(B,]RSG)^B2)C>0-6f#+(CTU=4E3>BOLg]Y/O,
Sfa^a]5(-D\ef>gGPW773abD3\:0=AdMM\M?;W,-gBVg9\D7L);9<1Kc?[fNOOK\
26/J5gI9HOaY.:+T\/g8>B33Oaa&X<JB(3VEHfV),BEF4-AGca1&K,ME:-(:SgbP
#1JEK:GVde<)=UL,DYWHRM?CeK4?R],BPEX0^=@=L8>+F.)gXDRbTOG@6U(Z<C9(
&\^,9UgR2E_]T^9[],/X1_ab.g_Uc\8&B1QR?[1>^=+\+d3[X1PFHaJaSQCE0)Od
AeB/6\[OT,g=cB<V>#0&L,1_CQc,];C(>Y7<?+FE43J7d5_KGe\WSNMKWL&29M>^
0D@<@7(>L,DY/K6R2:e>ZZHYc7)N&CEBH[KEK^N0fQBXLLT^DOa2aPAHQ@B>>Fa8
87dI[?-QT<Ib9G>R)AcJg>_;Z_L3H+;#?aR1BU2DP(e]OKA<,7\^b(2.2:T?g7e3
]eV_b6WfM,#V6?O<?LRN0_NR3>P:bXID0TDb;:AWOOGDbB+4EGf?)FefO]:fP&Sg
XS(J(:^gXDUdPJY[H<fI8W_-bVAT5E5FO8/,e\Z-S?d[a>eU9b,_:ZH,3\);D6bC
]]I_e2/SWHAQT8WaCFLgLL8F91^#aPDY0ZRWJUE.bGNJ6/f4+^4>NP-bYc,9#M5:
+8WQ1Xe[CG-=2>2?&_TC3+1&]VXD3?fJ3Md^M5bV2^GG&RUEB_\^/AO<eQN1>bR[
H#])F8N3dDUA&G?\E5-IMLfA2;DMSQfgLR,e03UYW+C;gaR1>IMZLY-4M)UdB=Ra
M..d.7,GM<f>feF^5I^.)OS\SL2U9[1BQG36Q#;AJ][C?AHCd6_AGSL3ULF)A4[D
KXSg?;V4&QWIKPJFXDcN=TY>dF7Fg>2fQb[dSP4g^/]9F0.JMTEN.,d8[CY\J]]M
df2AF8S1@f\=dYK-F(cRQC&c<;;<0b8H+e&:1V@0G29b[]Q?aEB6L_8F97AF-4+e
=<NVJ4KZ2#+BN1>b^S9P-3;9G&gP307cI_[<D:VHV)C:aQ/O^dG(JIA_)^Lb0VGB
I(&6)-bHKbH,7G//9M11e,9G3S0-1cJ6_dLG?Yd@=BJ9?9@Y6T:gV?YKXaU)Y(=)
8>KTAaW(\:YSPB;9\UF8LU:cIBgF6_eGGIN>389AG/Gf+?Ac[,+^OVeg,#@dUVB6
<g5=6+=B-GR2B[S9:?cIWQ]MGQG,QC1ZE7P@eTJB[.]cI6ST:M@@QEcTG;N\cVLZ
YZg>9O^,_ZGWd+FW3ON[?MTYV?d\DPe2.R?-B,=H1^BaPMEgSY7cQZ--P8QEF4:X
UJTCc()dA8](JP(#0c,@8.H[3P)SJ5b+d:.HH_FL7X2X#96-]=CYN-)?-^<]_^bg
JfQf3]7g[0eG.;95_d[gd_PWdC>HFeM&Y/AJ66cC=JFPZS8d=LR11&+7a@B<(Lb;
]=8bMLg(W65[^bS,ZK6dWBE&T9#1;FSAaE(7]I)<>LfQCRa5]^/^I/\bJ3&[JC;;
S:fL)_3ZB:2@Y#P&0^TFeICJC4#VU6<R)[(e^d:6Yd0_\&.NF1<6829R<9XJ.eP_
2@LQQ,:4Ke7AH0HKf/LZ\/fNQb<L=f7;4M&++T#g,GDS7(?>J5[@T/4JQHQ0AEbW
(^aBI;?c/+8<EH)BQ(A1^B+Zd6SW;MFHC+=:854Y?(1^ZI_[8+7CM;RD9ITX39b<
D85.:R34,da2)4DTPcR_;PREC?L&.;\HTZ(5&F83<]+4\9]1fe1#4L7IX0;?/R\a
R(9R.X6><W\[X5H2e7/aPdGc<-cF78TXa?/Z24)M&>#g<@&)NdP:#[AEHN)];a/M
F<ENM0#FM(@DSKJ1[Y)9-D2c2)11-,(\g)SBX/A3PK.3W2cY=)acXB^6Hf6c5>R7
1>&;LfXfL7OJ;9RR?_Q@CENR,(@bD_URbMDQ8,BE8aEY^G/Od_>1T/Q6UI:7,0>C
XWWT(E:3RAG@#O-10GUAUARO[-M12CRVZE77^,=F.#2;Y.W=M=X<7_\7U#V[YePE
cVNaG:YN0d9BJA43H7g=;SK@<EX[66\MM7.Lf?NU^<#f-X/3GbSU-;D<6c?)aB5?
)0O._;(dZ:fD,IJHMQEc-C]U+R-=gG1@_P6@51..0[GM9fL)E1]](SHG2YSd;M@J
F#VLH)Vf_T[S1[P<<6.dc)Y^MMc^;U3=?GZ(NH96_LTKC9:9U;E]QQb?,1VOU9RK
H^<gb2&<^IYJTSHQXG17#](NQGC0DRKbC3EO,H0CS+#>\M2ceA].0>6TZ8E@4Y]d
@fSR;9:\D/+?f><<&=H/KJQV?S9URQ]TaZeU2f\IfAH[Xg+5CGCO56X(K0O&LSH3
P9#7G=F6IHS?_QUTAHM-J>?R[J\C9XdD\.ff7IW4:Wd2]F[a:X=[NKLT,P;&fd>c
+<D6RRY?TQC,@UL9b&(aY;AX-J]5C3b>Y=#g=3)I,E4ZF0Ka\@bC.+A1&PQF>Dc#
ZPTOJ0acVS](>Lc8RE<Paf[ca7NU^cG5AG[Q4]8\:/)J&MLKKR=#24Vf?S0I,6gR
Y;;YVedVQ^Z@>g^:.[VWD?697UGbd(R[1SYe71OaK0f]U)LHT6FCXJ]=&@Wa922e
^7FIP\0U0)R;7?03aH<]RAMG>UWHbW,a7g;BK9MNScE870\XeaF,ab&Q3aecbW9D
E4V@NK?-aM2MFb-1bO/FWe>BZ55bS^(D]<1+W63VC^H@KJRYHa:VUR56\O.3.d)[
[/^P-F\aTO_bSB2,\d9/Z@SJY)KXg=6XUDK?9)DX1U\;#>K[4)eG64)+_6H8:Y_)
8DD9V.;\cF3b]HGVbCf>[/dU0=ca8,A&77@M/1R7S1NL>;+DR83R_ZDYKf(bb;GD
9a\I.MMR,>P6LcVC>#,dB,[^Q>OV?A3MI5B25,GGEG=b8+gb8:T,4MH1@^f@CSPL
\9[bBO=TOB_gZX&H2[dDa2?MDcEBaEdYb&+A:,FM7XaH5:b:2JBBNHGXcVaXeAR;
]<_g7R9#_cH;;T_@FaNFR;;<Ec0<T:be.6bI9_/,d+25VAN>,6_fT5LFSC]C;,;@
b2FBA/E=CZ(P2G0Q.c21Gc?>\[fHYBAI0&9Q7]]?L7W6=eeHW96bV?-6Y?R-2J4F
UM^:cKc^=VJ=FY;=:IJDD(IGfeVS?bVSgb&2AO^J)[>O>YgKI<5a\-VIK;^cHXP1
JZC))XZUK@[D72C.U68\d2K/G2G:96Kg\F6QO\95HCX7+CeL=-J1;ZW6\3HAgATf
B8OaP=K1.](BLad>-U>/ISBA8fI#]JB(g/3McLGaAY(d\>UH\DDWI\C=<FLCZ8MB
C2cA[JQBQUO9&P:]+.L<3XBSM6[LXCES.K63>(Xd(EEgfD,b<EOX_&X[YALdV73T
/N;N?T24:(7^V)d:B_WLROdBUI4H,=IPYYMB+e[K?_SbAEfZ(VF=U?#0Bd0I?I^I
_;8FB^_PL#ALcd&K^\SIK(VU)Z=^eTb)GRZ]POd?1>G_N0<>cGUZM\]g5f?56S[U
3>.F76SNX,Ic+YWb1Mb)=/c+ZI?)Aad(aLad#658IDAc9L+K(31PgQ@UQ;36X_Re
_Q->/WD>ZI;@[Q#AV^5?_JG41WJ?R]Fd35f84SZ,G0fJ+PK@Q:4bU)4-]/_=1;Md
06(,#\#:MQ,,aP7&W^X8DIJ,:2HGZdN6Oa&C0^P]J=[>^[SRBV)L:/)2d^@[G<+(
MU(R>-5aQ=]2[b02aW@\UV:/W]\:5)d8Z(2A1+463ZeWE86)695=EKTM^5N=1Tb;
YW\\6&RYVb_O6:EAcSHB5[F2@U&4WYT64X3CZK)9BRbCU^5LP?(XfR.0DGRHcgY^
eC#f3YTg+a]d#.D)/&4W@5IJ=NaJ]9#8IeG0>--LMZ4#S2M_C:R5=]/&<(G:;SI=
31XW<cO&=5[SAEZcGXW4a65efU5F0FTI(aO\P(WNG=2fVSD?1.S0=@Z<QYd5#P4K
_.1VD<.7Y8=cT/\U^P;H&^_g#)[D9K\H(Z^Cbg:d8?OTIU./])CDFX\?(+FT8-&P
?C18LY;F+O3(VS?/_^g(R_?_I<I=4X1a7K+cD08>#X821\(.P@d\A(L3,c,^&g:Y
W?bdKC51g&f-eV[Dba&OE2D@CFY@L;/Y@Y\a);?6,&=-<\K:X>=0a-:b.QWGFGa?
T[<W>/[UE6QD^-9Wc8?UBM?/JUK2L7X[-IFZ+]e@f-O&Gg\D(M>A_gYbE0KeJK70
^LDfIU]fP.V=++.A#25Lf9\LZ+gf]KC3/8Ve([UG,SH:c#CI&@C<;-[+f2:Z)Q<_
9&B\A3T,F=2>;2@^GgD<\F.#>NI6g\USIN=,N]gd&ML9;G3+^aF(abDURK@_W,f[
.2^TO8,(91RE4X1X8)QUWQI(0\M0-,bBU)-IfV)IKC#[.A=+3F3bYG9ZJ[RT96/a
T)+cMF-egefGZe/FG7Ub>Uec+-4MNY+Ja.-4&AVQ@#=>OAZ:cTW#-HF[M=6HCL<R
EW@_IMX300LILa6]8ULba9,BCW[#O;LA(YO>C4da5E<S>??Q+;(E2S0X[K9CSXIG
fV]:YB:SO.QU+\I.@Vg@:2C#B+<9&<.IEX81AH:GL8NQBLUT:1=4Q<K@&B^.X8>e
(+Zb&f0QL2aI=^L)HJ[>/P_BXd7YY-,QE?<_@.e_1SE+SF2,W],a[#dMU9V>MN6Q
B@5O+dfQ(5KKO55):P+47Jb+0]QET_[SL@g4G[J5Wb#=8TL>J392eYf;EB^cK^V9
-XE/65Z7E[B\a@-DB.f+#B0_E8I<cS4Fdc__\,,,VLMU_aBW\,EEdT:4SA3E&_,_
DBRS89:V_c;:L+4[dWFeP7b4=+4)B^-J.Id:@>1DW?aY6+d+ee@#bT(><V=+YcSF
C^R=5,KHB?2?8U]=S[2S^,@J>09KY).a_]WG475?(g+/@g<f3Y.BJA&Nb<8)-2F+
^D8,P#=3@5=3<RD@C1F)SeDU\],J/N#.[[\F5A>(eIZ+R#QHNBV-@4[8B?W,fSM]
[>\_KZ)ZC9@/JLG#J>A8DHG;?gIEJ_XR[44:ZH;QL_DFM7dHUP,-F.=5&8PQaJAM
[2Eb.#^<@QD50R8K.M<6\(Z]:13G._f@>R=>WBT4X94\;_INTT)13G6&TM20CN4P
GJ&7#D?.4+@6NB7Y_[76PD[G1M^YU:S2FfG[2?EFW>HeX9)fOGg>A(DTa/dMJ8(c
:9S+b>:\<[B&+4CKcI^7_/5\cN1I)G(UKQ^KE9PDbcWO>(5F^/L:=e:T27AQe2\d
G2^3DH;>+?;IWfcC-D@.EV.f<Pd/62:g#O&&)^\e3dB8TIV(6dfR#XD<5=6GgMH5
74g8/1Oe\(]JG.O[=B>IU1ZL,gUY@K75.D8T^5&NI5HJ+b,OPcWf]],8K@HX0DXD
Y4MOFM18g9f<G(X?58@2E(:b;f4NW&^1HT/3B3/-17@K:bKM&//05g];&a7B7,9F
HJDd1H=#AB<[DF2?T6Z7]0E(F3=/ffgg^H_8>3?I/8+6H1ga;-eY<G^+;H82d(82
#b9g/#X@X+7XKCfK7I)B]N211D+/B_OYUY+c8\X749b\53&#<CX>Z[/b=/OEK#FM
bG@^&^2X]&RC+J+TBE5cZ5a59828U5@L=2-;H]5Y,A0->B1/)bgB2ZCL/SR>O#JH
2(DDI8DD9gBR:<R(gK?/e#T8EZE<0Mb8DFYaFaDUAIS&?8)dc&@HBL>bPQ_:.+aW
U4:)>cL7@>AGL-Q0A+E,CeeZ>R&<K(=I@+Cg-D&;O,3[4()2?:)I\^0P-#/G3GBE
B1+ZDM1\X1B7J^CO-;_fTYO4NCQ#QUO0FY#@3V96)-Ee(B2L1,C&e:#5@Wg3QW;d
e8>K87OJL9N-50KLf#LXb:ecW;C-KH&_VN04Q0TPOP]7C8\4\7@F2:gRR7J8dEF=
R-f083?1#@4M&E:6g>CC[O_;3bA(E?@H<T1-P7L^?J#L.6-bRNf;2OX]6T][c#>Y
?F,=>Le0B7@4g882/+d6XTW<GG^1-7?=U;9dd2=6c2L(=Z#3e(0Sd3]?edQQ\@)[
aAVG.PZP=:&Bd8C:;gZ(gW#dS,0:OG^1FKM@[gaB=a1+)N[NWeNRd]5O5Q_-5c>K
->64aceX])Rd72)PMYc&IM]cZddXC@63I9Vf^^ME(GV-#MZ?-NcWAA7dK3@Y2J>]
g\16NVd2Sb)HQ-YbaW]C],:Q[M(GC:<H.4Fa&OU@CLJ3EC7OE1GE6UC3B_=O4b&b
TG]<_;)M91?;V?+061GE_CZ:696A/]:N>#O55UW,UZM0(2bKa?3&c@^\,eD+:7U.
-7G9IYN(WfD>G[_X)L@@F--Tg:E4T]()YO99B7G1TL;<B##)VD)EW4GR[N1(f?aX
P)FCVf>)bUHT/_gNg4F<NEKG#C9Q2JcGdHCM-\DEc1eT=51YS@bS0g>[GcGNg:-.
OE?Eb]ZH^#4.WGfI>2=_XG+b@XX@A_SVaY#X@IQ1ZJ,S@\FN7D>(:>-<OB3Q]TV:
g-F-_.>VfQD@b(+KJEL7ROEc&L.)Sb_K&T>,_FSPD]TcN[()M7W_Y:XXO@6LR[V+
[d=#0@>?85R)M\EYZ:MfF\QTd&#cYgWMOd(_:Ie)<-QS3?2eP#_7S1,dKPGXRN58
/34IZ&@1PIDf,^2@(ZKeI(/Q;QQf-SFMD^>OecZI-_SDR5dWa[VL7^+LaI],/TR3
+^+ZE<@I_f;d6C?=d06SX?LR&/)Ed.gK/<&6X)3(D?>/.29MPL\Z1&=P2#_0<3B0
];6fd5d13g1P=0_XAUZa5A)_(CAf7)e=dA.HUTC8G7If7gZ&5+_g4(e1N6d^Q2,5
EJY.[HbVQB/#XLW<bX1@5,#31S500^0P)fDEfdD;=>)XE+]GSO#05<ddIf]-[OW8
a+6=X/W3E&M3.=cO3+ZM/\b@-44C(N;=+S7.V.#TI+gTM/N].9_G93F7KNYDE#:A
Rfe#H:4HIXO&O1AEUN)[MUAgg<0^1QWM<1-_>eO,&=Qg]DE[[6E;Lg_b.7[)e>^<
,VZ/@->g+f6#/&^T@?+Z+SV362,3IELPQ?J=)e^K43J63EE0(L41D>;CY@>G0\77
X;[P/]W_7^2-\Wd>Xa<YgGGIO)QR#e39=aH[=85dZ:KHG)])eJd26c;35KT)6TRN
(W7)<gVe2]LW/fcX:D\GSA+Z(@WUL.A95ZE_XY9WP_.#DM,aB>_=SK+PR33ER,?+
=4E=NTI&&,>IIV:eE\13f<<L3.FEG9fPUX^74N#7GZXKaA]YYD\MWH-K#)HW)XJ^
KIH>:Qg1OSEg,E]JQF#MTHE7V2C1BF_)dL9V3/CR&P3C),:#9ZWfO&bc,^@1\-67
;\_+T>c5Ua@UBd4dZ[^8)J&g^FFPP?DN14@fY4R>+:ce8^T/?#39?H6]901880?J
6_L/U:+<=4P0-2//S_RX5,8MR_.FIdR_Y2]_g2cCeWTEF2WH]SJR:S,JD+&ZTbLS
0@7[#ScbdTRXS>b:BC;@DDdc:OWe9O7&Bf4[:2f+,+9EDR;\eXTS#VD-g@?IKZ?W
X<:9fTgfV4PMO)D8K,B^.#I,BFLJ6gHAAa&&[Ye+UfUIc[HacB(a6<_,BfP(F5]+
4A,JTeSS-eg>V\+K2).1H64cbZHA>4X0]DcD/E:&)BJTI>VIbac_d;B/PP<4/SRV
6KXQF<_0Ec^f^d[,a?(O0\7f_UFSVA?#=1F4XAO3?fCQG&a#E:1[CgC8J7gEbM<_
APTSSRJTQJ4]MHR[S/>?P?>(W]\AgM@#9<VAC6?[EO7./Pb279]<>ZA/IY164HQ]
4E[.<&b\O/(gY]2g-I5S&b&X-G&.VZadA9Z1d9FP<@OaIP+PG37/MA2ZE5]Z+cSc
4,AL5=ZLeV8JFCVd5OU-.+8XLbH.c:-T<b-M@M0(RUNWTP;A^f_/C1/^XGZgDF-=
IDK717C4TIUW][-Q;STQ/d4T\(/:0WS_(T8fG_PCL_]Ac&cW2T,e^RBE7b+\gFPf
Qf@Da4.eO]gNGE&L:AGFV\)eU:[4Pa0G/Qe?fTIPYZ88].J>Kc\eB\.BV)a>\J:;
K#?<XKEB272ZJ;ZDV-M/G(LMbY-OE@-RLI\C-)=e1D.QRM/K6e_W:,bZZ0JP/Fb.
.80FRQV8&J\P3fHR0c(eAY0gLQfPI]-J787/4;>8G12&9K[FXD?626]EcF#LJJMC
>6)Sbcg#L9?JUFY:3N/U@T]IY;+X15Zc8@<,)c0&W;#@23>NXZbC2@[cE(eFOG?O
32UTE^W\c=-B6(EW;27[9\]LYXOY3_KJJa+L2baRE5[XeL5@TX,/7KgL1K<Be[1J
YdNOba.\A38a5G,&)7g67NKYV+=FG-4,b<8#Y((\@0UY]b)I7?PbI/7L31K5N74)
^K#CfH)#TI4,^FJR31ZV^>SL((#/1W5U<W_;JO^B?#M4(O69>./HWD-AcT/fON:2
++]=&ac9:HI6O.Z6Y07fZgJ9;]Yd7582-@JQ^a7g2)J,@?42N2J<VVI?=#V[[a3=
YF:If9<,JR^YYTL?C,DC&04>/c>G<X,+[H#39AST5:54P^+N6\?DF(4J/ET=dDa>
BCXc+F^G]\f?Y2ZLF_3d05c#_R>(/Q<f_gN:d7X-C<[OcZ:P@NQMIR^[gBdC8AKZ
T/VYKSE(/24fK7HF/WT7--a-.0R&ce@\9TZfX)[Q>R;BQ@OQ.:XQ(R>&##-M;;3-
IS8Q-Y1&SV/b8W=VI)ac@W^8I&4)\/]?=E]][=?/O/ELF.dZ\7ELK:R^7SD^XE5Y
3aKBg40X40GBYfgS;,;04\46ZU?&&IWYY31^_6X;3MbV@KJU=E=f#)Qcf9&?BLZe
DbBC#D2=,fRYKPU8+a1KT1A-UIaE(D2F2CU@?_X231HBL\6L-M:/8^Q[L6A)=_Y>
G>A,-,+G2WHaIIfHgPI?1R>XS:V>KdP+ILAEX?RbW7[(0R,c1cRLO:dC7GfgD0\4
7EO+/=K4WBX@)3B?U44OP5Oc7N=K?K,,&>aSM?=6c\/:BP,F&<C9T_4KeEGE8G&1
,8Y/SDQ2I/)RN7N.PK9FH[Q#eDa>e6HPBg&OOT_(C#\2Ma\R7).Me0VGYg0B1CO.
2Q<RdfNg-aa\F:5\V9Fc/g)<\/>LJ35//:/MVX>[CD+PF=H>FDVYeZG+OVQ^?Ja\
\I6SWF(I@b_M7K(UaKV)Z=\DA3Z?=S\gU/S:XWf/QL?M-B#M#SGaV^WIf9Gg>[Mg
\cecX9fNJCX^\^2<Md.U/829a1DO7a&S7/)NcPDRMX19(^CTGW,YAALWbBS4D:)T
VOe)(/WUQ(@g2aB+cb0AI=(Jfag29B3R?]WD[Z:EGIGc-1fc;T#,/5&2Ed4-J/[e
?P7PI_<#R_I<NSI]<_L6<EHY-)QW3>C=+<(GEV;8=bG\_2_YM_[US+3?/)V@C-X6
,L83,5+-X;1C2=S0(&)6:2K<-1SgS>#ZJ?.aR_c)PV3XKXgYVX?I1.OTJT>afJ;-
&V;b5U,P35.<]CQdFY;&(BQ<S&EI@VZWHFS/A=[K2Cc?6M1>/IM07;6E)M0QI31Q
;\\ZWgDP0HINT3S/BICF8(<6EN]J^N6fMWE-S>H)#<[_T\L?DaDE^e&fM7</UL9(
^USHRMNg^5Z_TE9b:M=]aM+:O&/(U?[TL<W^40abJAJcWM^\Y?8DaL.afeE=Q[M?
DXF_9:d0MG0]7+/^=B401;:\]G@,\+NQ5#>6U^V#XV_@B_I;d;a[Wc[J;]dRM&+Z
W)7#9fW(:fF3HP>f:U_9U+5a=-c7L#-WBDWS(2eaGGZ)FP_1F2QQP.g].X<M52PJ
8:5(N@\]_&]M[\\8UG@[JC7KWSU&XSTXNL@3bedN6G/ICNGJ1Y[TNZD@;3DL@++]
F^&VLaJ0:DB2J7/+#</>041;f)(JC&bcJ[;LdBLYPTV0SS?##-/EaQ>0<C;Ng^:f
M1)=WXL:,V=#<I=:5U;&\_\+<d>6MgOVcGNNNK4NO:SX[cA+P<=GS45J4?gLC-],
UHG_=77_&G76C,8S\K)O-g^(&76dZTD17CD+d/2EFA3^=ZW(QY&=4bJYU(]e^Q+E
Y[-7X(];3=B-(Z@;WX]N>[FP;3\\eC,06?/TA7Y-;J7[^cfH5/3DgVL?g3_E.a2R
5-GS_9e7_;Sa]ML1FeJ9]gZHfbP]7KV9ZETRP4,;5c#HKVEDG]\=O5ZbPIN:XU(>
8f^\+b0dPPZ7ZQdIcfGc5-Og9,A_N]N57D[RJge41cL;N,DR5Qd^MUAJI#9/KP7M
H4V[;[b8SUNXbQ?VW]FJ5AYP-TE_=>3]Q:,)G(K?8^1523Q=)\)FF:V/3bPeA&?Z
-BU50E?;(YGcJe&02d1Y/U+g_GGX<c-Q;UfT6+b\d<;YbTW92+G2USIE>[c<]6_d
>3U>>b>1W>25]R/YLFdZG25IH[Qb(Y,H&TZVCUU+8;aF4-a7XBJB(]/Y=EW-I:7;
cF7daDYP)L3_H\HMF2/^9HZbH/(?8BOAEc9agA(XRZ?YF^5:]ZVV>(VAM5-U\YZT
Ig=6Hd#aI\675DbQJ.>H-+VAZHegMdfHa:cVeTT,+)0VGc-/L]A&c>9E7O7Q[T-:
J1O,LdZ&fd##=[D^<0cT2T50>B2\\KXB&D+c>8_EE8-a95I?)gOM/#bZV;MS-.Hb
U2_H;YL_GIQHSe\7))8Ia,/:c\?9PO)#?.6#Q[(UYNM+#8K=5OA8187P:=^aMD<f
L\+B&X+QLW0\LW79@O_+(R<7^[/GfPF7_Q5Fa&8A8AAWSa0-;;N?T#6WGZ8-ES\N
JI]Pd?J<+<X9b20T\.J:)9ME6gB>;0;M2c(^>bX9]6K(+9-0#]QDM)13TLQ/9Q/6
X+6GdcBLWO()L6)1381ZZ712Q55gfMG3bBTDHL_bDU)Z:KJ(@M?1g^.@S>F=F^f&
D8a[;EbWQ-;##S49XX[bREIX5fJ:Q;NFaGS_??G\cQBW_V,^>7>d3IYX@TWUbI^;
?<1&&cPbE=RE6[:HMMWc2=.0eX;39V6?g.84d<3S^M8^J()a:#_9-Y_QF[L#]NIO
,d#Y)TC\ET.Rf\KOMg@;P:T0Y=NYUN+3S,__VVgA?L>J]A;.NKG_GTM9T)WZW)gG
BIaVVBURF;6NM,QSR38^^;AEASS#TNQQX+]4,5=-U9^/(@2M>]5R1gf?:M@PPgBD
7?QKSYEdLgBA3gT?-Ge]I5)cgOX.VE/N?geS1aU02MZ\^664_b\BN&=AMEWB\\=I
201OZHF@<8<-&-8;e29fFMY@8A@NK[I&GK]A;N]@R46]C\_=K@3_S6b3bP/g.1W.
/,M@Z543HY7,&L6dJ=7H]>6\,=UM43L-TF^=/OL?Ee0C_3e3Q[[BBKV2PO[Ca:SJ
/M)H28Lb/D@3T8TZ,b&9-;J3WbKYBNKOBI&\bB,#:c5L3OOc^?7Z[(YXG4JWZe?4
N.O5E6-[#C^2VAX9VYgREX63[gN+25&E4<dXZQX#g640+G/ON7D1P35RgBgd=__8
;\NaP:BeY^M\]#2._9)-=V56#-8/gUBP?R05J&-T6e8_JH9#<SEO)1BR-T\08UHS
8)ZTg(5ge_Gc0E8\E;BVLZR.IWX6:bH3Y4a/2K,HV.D,dRdR?BAY2Y^dJ@OLCW[M
IObX.,/L0,M0T]./Q3ZBYWM:gA3MVcc4#P.8RK^=XHf>]AY?3U;CD+?_VaLY^GeD
8/A:,S;,56)O,HeJZcRP0;M?5FG27M5c3Z-TJ#gFJP=_+\6Qb?6d./_g:EW25=Y+
NBG6Z]SXBVSe<2NZ>Q9+GHJKcF\,9F2#Ob1IW.J+W:X\:-:&G-ALdC94;gU0H\W#
2>A;Vc>>C1a,VE[BWNDO@AMW5\M5YIG7C^e:VWWeG]I/9K9OBV[a)f6AOgcH5M8e
H8D=23+>YafB.NaU(RH\.@-gc_eI8?B5e7a0H54g^NGB_<QaEgZIS3ML4Gg]-9>)
N6-VTLDT?/&7B8.QD^.6CBf>C/cB?F+BO.VVc.;@:Q,#HD=I>T+(X^1)eJC4/S^1
g&ZbLO&XT4#WI.b[8B/=XY64bYJ)PFAdR1T7\D?6a:/9,0,?cF9MP./0]^HSCH[0
LdeQ^QLIOL?\0ED\TNWAM^N0Ed9\=N[,Y0Q2[L-\&B33<a]BA[>>_\>W^68E[@Xf
_H2=U/M5?82Of58;5/^2WPRKJ7/D;3\-K+_50Uf=HaNG4HE(La#5[O3VBKOP&_N,
1G&5\.25+a>H(dSFCQ_DG+I:FJ0c16723.0.<Mb4\a#9-MI[-KF/D,3@2(.BNPOU
2+e=0.Bg@/D&EfRKC\gZ_gc2Ld)@Q(4:^S5aEB:;2:Rb9K^^fC:#(JG8U/>DECBK
f;EOL5Ma7YBL\?I,,(TOPN<4RKc(bWH09P^-:\IN2H[\[XOa1U4M8H#P^KR&BKM=
0MG(9[9AfTbFG@38&.d8M=H-:,DQcgT73W[M.^X)UcF&:=:V:>/W6NT+^,N+YR7J
:<_YLZ(U8LgVGT(6M1BX^81^FX/2G_4ZABT\^8Qd;O.4QV->AEK&@3?dSH6;e5ed
S7PN)FX&Q1g0<+N1=0?FLR@T?_f:56^F^c0XX^Z=?.@T15I)b?YIg:+O&Ad24ALX
ZQ^Ea&@33=9<T0FTD\8XE9AAdcJ^.20/bI-.F^,6=S)B;YO,C?Y5d5g.[Y]0B@DB
^fdWMU&9L::QfAGN(A6)4M4W14Q3D)U5Hb4cWX3,d@bR(Y>3_\>ACBV+-;,V]W<M
1V5.Ge^W=g^?9N^8WVF=K9>AW[XQWdPgee8R..YV&829JFOD,BC4W=\=F;T3bEQb
BY0dD06T?Z)TWfZ52YEI&g?IHGT@2e&VgE@6;&3a079A;<W-@WQM[GH01;TXOJ:g
7PCYV+Y\W/GTP1:Ib\X9GS@Pa)\e\bJK6I2SBS5#eDY;<BT?\LW0_]?]a5#]c98C
U(<J2Y_e9R.,,2g>cPaC2_]M8LHE2S#->43E&OTZ[a<^TZ7;gNOE[B+K4/aQPGL)
M@/MUIPVU];G]MMBg?YTQZ5\UD_E#(I2gZHR:)J0Dcd55#LTa#fd?f^=Z3<MGRYP
&4M)ec=b?,KT8(E78L;]I]YI+^W.NX::HY@.)L=/=50.cfWGa=+V+g>S#bE#9Ea(
2@0Q>Y@RP)AN-f7ZK1S1+9+@TO/H,Q1(P]075^(8b&f@[,?8KDT;CQUg-S2a05H>
<AMB9DF0\gM^^4e8+]34SDO,O9;fZKF38W&fA-UQN<g.U@dDQLMaMP>+<:Ha)43Y
2cN.Y&Q33?,4/20+fgX9&(W#A@]U[[AEe&-G(gA8(KfNZG?H483M/_])B\:+/:dc
JB\LVY7^ETX4(Ob<5.,YAXY+aB-&A<LXZMBA#XNB);eES^)gO,ALbcT\I;gQSdI@
<Qc.J3eR.eI/U&:9bAc^Je\f\ce=M7>O/BM0D?Q8Z/=V(c-4@T=L1fXFSG;bg#)_
Z)M.Cg;(MP[10bJ(W-8R9_[C&ANXC=(K^HE&Od9\?I)^b;8.O@J<MQ1SQA-GIfe6
<ISQKSY?&0615&06X?^?;PQ.>N0^#^?9^bZFVc66d\:01/JGDGWeXN&?;c4LX1(_
CZK5V?7;>_Hcd;f,FH(>VIf)S/,CgV2EYPD5@QgM<V)L<gB:W\Z5g+C]:HOC3gHA
I6Kc^_fA7?eX0ReS=9.I0VNT3E:TG&)a7-9_=Z,QZ6K-&C#H_Q@bP23?LNI+c=b,
HZDAB03CTO;fGYFO4T;(:7ZOAAd##3F_@(,JN0>eLYKRgeI=]YGe@EDGS&993JJ9
fa([E.R]/ZYNDOQIdQKTOR(;9SIG=R&TD>8F54cJ-KF&8GDBVaNC:D^?WQfV&3Pb
9.V._&bEOWC,=AUIa)Z+9.A.]#]#;,[;)H]T^KcN7+,K=f+S<3OW]KUcVM=EcffI
V=\BL\?[CXSH0?Y2]_L@O&GPg=]LB,_9Y,]2_4,0[f.Z(2(SG:6W#\Q=G6QcMEFT
/-C#0,SX7E-2(R7bU/A[1[0#PBcJ]GVN.d7;.:NAUC^6(3=HUfg/C2,7E(MO:.a[
)9[+?2:+=XS7ZFAAg6V[_;Ud9]Lf+WC?<4@D>8I#KIbL7?b6#3SbE\aQNC+879WB
SO^]3aSbR6HD^M+2)@FB).ZN_eTOA8F=/)WP9?_5-Z)H>,5&J:cHB<Y,@.S1JY?E
S&_>7XED,G&[^6-gNX@L):^AS&FCKaY.N;-J]F1D?ZNb[5U4dDIJY7^Ug1b7U?DV
caaE2O=V[E2;?[X8</(ND._6HC3S2Z(5Z@Oe(?XJf@Uef-7,UebP4Ob0.DA/XFcZ
+5:?,3,28750JQR+#H_/#U9TLJS:KYPeb-_VcAKAAVaJ+C^8,NS4:ESfd4).47a:
OSJWZ?QV3.M=YVaB]6RbMR4/T)HSY_EBNIYf.@:/fOS(-E[D#^HW<JWg\A/ATdFG
RVGL6cYZV\fA9XB,\gb.8SVdOFa],P=+=JB[\)ZFRQO33fHO2bI@/I(/+eU5eS.X
BcZgU0\D&7\O:9)H7XJgAfP>[2aCe,M4#6fT-?#6Rg.4&eZfYUJ)0/HVKf81@)B;
:=B_I,(XEZ5RFb=@S09/RGR3G+dKZ><LOYO>0G(TBUX(EV\)Q[)?RfS7GIc,IC21
=O]b#L&Z+A?11d5C<S2.MWa;1@M^>UVVYKV8[HbEP&]GaFdI0&fE\8FRdRJZJ,9E
d\.56GOcaZaC7=/ZHKW5&/1bb:^d&f3,7:[XR.(ER7R?K9BLX/,6JUPd;A/f0&>5
GLRN7\R(b?N0AW-S99fT\g(G1NR7T.98b3>_;07?>]LS#>(7Yc#Ge]O^(9e;8\RQ
TONd&ODa,Q+5/=@98(eL/<4)]48d_7NAAM[D1H6\@:AAbH5#J8fQRA#E)KHW-cbg
()af.A-Z-3\1A-HVIU#20\W3T\.)3XfZ-U])8IU\)[g35OU5DJGWd]bC(I0;b<MZ
E[a8cf0K_0P<[DOeT3?^=+Y,eMfS@[c3YA5KI&P1LX]OHd_B3[Q6N^Ba;BD^Sae5
#HD2]0f(,TOT;d:SLD>>1))DZ0ES5)XVR-K2H(TSPKXP_E[M#67YR0aeX5E]U8T+
+)AR/CDP:MT>]Y<BGT\G8,gC/ZeAXO@bLSR7/N>&Z\XOKZ_4)G@R6.S11_#-#e0[
e>RS/aE5b9L7]E1#NTIf7SG=MbcMM?)9[IE;;[X?ba+EK:ZDHc.A<NYD[9MDV_P1
5>6;MG0KH4\HTa50:0:TMA#5GF/;cOS;+ddBP&Nbdcd=2+#Pf\\6N;JAK+9(Te<>
0dR.:PE0H;H&)_^bTS]#OFKS,OWBd[+8+M8f#;:If55+M5;YPgeV.e1WY1KLVM2,
Db^&bNU^;W,+&+.dgTE;6@XY,):I6c<Wb)0[L>;=,3=gZ@f.^OYL(47A5a@bX\#Z
JF3+WZ]aR#T\EHIJ42Y)d+3]255@f9.e,cHBS9W8,&bP.O4Ce,[,Cb_D-\]V^IO_
-GE/MF];HXbWVXDLQ^3CBCS<8H><QA8JC3HaL5))c#J9^-8H3+RJgD.W5+,Db[Nc
d+??#B(TJ/aH&,Nb,Ue5B?:,6E6A_cCR&)=+[6X1_.P(I_6>^@VJAaW;+OQU?+,P
f\<ePXM+J4(<\O)S5,eDO>Fe5,4L+e-bQK2XF]Z&#A#bg__1;YXKbSJPeZDS#]&R
4fdN-+P>72/(eL#D3^DBKJ\QG#=-S(OEST4BbXP(,_4d1^U@aXJ:PbZ=;\BB4HgY
0d+.27^0OQ5G+>W;<f/&<fJ:@7/e3989MfN245-LLeR>#B(I\YRJ;&,>S/dS8Pg<
>Ye3B66AG;Q/BPTCVNQa<?Yd_1Wge4U9.Z>;6K1X9aTZYGYB1,G0b]fO=bPfb_75
HXT?R?&eTO2KWH,_7=KS<(&C1H,L@DF1ZOd0X_2Z0V8G8WDY#:^+RO6,/SeR1FUB
Q(C\J.=RaX1B[=F++BZ@<VGPb7ICJ,)(f7AP1MRRcGC2ZL(PV;dLV=a2/.=6+fg/
2?]J]<T4e>>P7&+Q8g:I=eUPP&63R/RT)D:66ONC)BD->F\L3WKL68:):(f1dW.0
+FNBOGD](2NK08cX&9(@0]=4J<<F)QT39W&C:7ZTbOSCE3L]<9L]S,P;A1;^dRGU
Q9\YY=]9#1=@f=bA?I-Uf-;HcPS9WZ^8EN[9aB@V#\>0FeXPXLI#@a+a8[]A5=OF
c-Cg.1OC50ZggcGLKI8HTL\1TYP17;/E71+J.91X^4aM/A:H)./,HA1HQ\H011_g
7A7;VH9S6&8g0>IdD/&@dg;O]9+G9b.55>Qd>\[2]Sf6gM136dIbg1+Kd4gE?05S
3^Q2Yb8cES[27&RXK;=--ZH.gA<Z=\90PNHO0GbeV[D4<c[fET6OW@[E;SIHTM>8
0Wb832,OCdCg4f_GF>Oe_@5b?W+Rg6VL\bAc<cOMeJN4-R/4)NAaSIIWPLA0=#@#
1aU;WFCOV@?\K0XGU<..LTFL)=7M.:A;=A)[aD5)4)(.C8BDUDZY]_.C3RR4&K]+
J]N<7C(Rb;8]AH>6C58C-E8d+SZ//<aHNE(d4:;WPbNQ,ISQO<8Bf,AOebE0M(BN
[2d^HATYe-f.bB[)]]a3bLBSb<^.OfH:Y=WJ=0-BZd]KKUP.:3\.HFUA)[NdH()@
RVLe:(D;5aeBPgb/4DI5>dXeHQa5.W)^H6eda0]fUZ+/R<Y.O.8Y#?S^KC4R<G]8
L:[YU)5>^cZg=c@RL_ZK7:@deETJN)0H,;ag\E2;2bJ_,1\7&/_OX#ZfI62VGLdK
(2>Ic@PeR;JP=U8CE/PJ+RDDb=c,89L>&;dVMLEY[VH_P441E+df=S1(FPK]]J4a
L.-1/QIA+P^22=[R(eR0U-Ke><VT,bE(7XeXOeXE;be.=8[>70\:;\3MYV4edR=d
/P6@L-S28CbD?Y=@)01P8]>@?OGcKd<CAR4PHSdD5)Sdb1)F2AbXM;2b48(XF9,L
:DEKg-3a_QU)RQ<e;Q]AYfA#\aMW&E0QbdGF;W6)^Q4@cBAVTOb=(Z++#eY+()8e
N2SYFT#GO7E&581a=N#A9WU\d8>.EF@^#/DB##N=Q1f.VE&GK]Z10ABQ79]T8Y^_
G)@<b7OZ<6cM=.>\FMU<0Q<1e]U,:BA/+?@8[dV-P9E4;c-6T_,GcCKQ7^,DD65Y
[c-Wc73;@=]ZET)S8YL5&IN26_UK^T>I39K@T_]JJLW3+6._&(S+MO#CG_)eLV/X
7:WdK<Y@,ZVWGXcT3I>@\)c7L(Ca-TPgfgQNePU,=6ZL@Y+e:G7_QY2G6dUO.2VU
HP[/E^_DPS/I4SFSLAW\a2&25_O7/G=gK&F=RBa0WfXY&,_[^;#@a(:#gDJHE(0H
d^S6]dU)b8UOA_1^5DV#3^Q>S-Ufc&N2(@Rcg(Daa<L/>EQ^5agK=L)>LVX.]dH/
7WR4bY#aB+Y0384BOP^3.(MVbT-&/PS]PN4@U6I]6F]QbD)JO63[--[,T2_EaXYQ
Y[I><,4Y@7>Z:SAR9IH7P/7K8OTD6WeV:XYF<F5b>^eYQcPWG60((GdGc/Cdfc=)
&:#L#5NeABN5Y+TGP3#QdcZ4EgcZA.>.T##NC1>7d-OW5+Q+19LV-QZ;fO^XNTT0
V^(>ZJI_=]#U^abJDNRf/5@L97/CD6NEGHa4P8<0]gQXH#Ma)bE(IW3)=<WdS[8B
8MUA[:6]^Fd/RTV2]dg),QI7gZO;SL2Sc5;MaBGX^dfVZTE9c2O?\0)GF65LEZ60
S.OC9Ld5Fd;66EObE\=WX\-&U=8(XIQXGHVIP_DGLHbE-Ie.AF9e\ca_6:^\1.>7
AXOd/F2)^)QKbX3T9&SaZ&4D;@&;7KZ?]LX.Ub37KO_:&,_]dQOReg(I/d5(-/d<
@UU@^<E;FGPR0))dP2^gBTCMdO7Mfgd_d2UY>LF=KK+@8K,T^FSfY<E@H]PR\YVA
b#VS=3cVe<\]EC?G&6A[+=f+a1f2SV&^gPfPg,^C7Ia^AMY:4T5g8R+\:c,IL#He
2ODE:0;:3M,CLS+.\O=]A8\WXGDf[\bBNe1f2901X,8^3/#Z+^54^K0147^4>AXQ
T(c/^6K1=U:FO,ec_DRgJD,2;/+-H46g:a0eLB?.(f)W7La?<(_8;DSeHG@RJ+cN
(PS=29d;B86,P=@LTg:A]G]\,B3cOYd2#(Jd@-X.T.PQ]I8,HdHX/VRENAFLSFb)
9OP[^.X:@54_Q-,=DY>L[.0&P<[9=6]5H@]+ac=Z1]faN6OHEa[CS_]MdYgMAGgY
3:95E2O+Z/0/E^X0bJ4G:KR/=VbG>4:MH=8Wb:B7S#g>:;N#MWN37MQ?@FSdB]+Z
a7YO-+)&FUW+BBe&?1_#PeM2QN/9OfV_LB0(gY2cG\S?73RM)[g[YWM\G469Y1-S
,dbC0:<0ZTgb4XL;4KOBb9AIeMEP6/e;)#TPg8Z[5+_&S>32.OZUWO8>Z99e1Ibc
.XAS:eN(.V;+TEVZ=_=^eD,-=/fG8-M0>)9\f<:KW,-4O/7^X\3()(9(DT60-00_
P?D-aB6T>1AZGG2W4O=8ZSLb#3SFF>;L[(6cWLB_f6/&/C3;fa<B(](Z492Fefb8
bLH86S3EATMQ/QB4\8@K+cf#ZA(G)V+0<06A,OJGZZ+H.,@:,Q_\bEMQU@ZEEC@7
3Db\6AQJf=IOJYL>e6[a7P:cMDF^d]C8^Z+Ob4=6-/W<QAaDWT=ed]^FdRLJgH_Q
c#+ZMPGc8W[eV1f9TgG],\J\Re7ag(<<S(Y#U_Z,Hb)[ZB-]&:P1b0B:d\4D9CYK
V0fI+O^cQAS;XLe&6?@:-^/WdZdEOLUd1\_&Y_O1H3P;Z5U\^fJLK?@7:D,0(0N#
PVB0D7BK_PR0)O-V+9&^-F/QD@TfZ]W;U[XIAe?e,9X((QT=3?))aZB2)@XN+3P]
=?\gZbK?T8;3J4a\dMcW1&;PK3O<L0fGRUDD-TK,D^R_@RHO&d>O/G-C5O4<AK;\
_dQSCAY7<AL&U6XRVS\S(gfBQT9NMdD0@M1:A7N7DcJ&CG\&3@\/b:B=d&-O?F]F
ZJbDDeT).&<[=/a&Rc6Z)7=9b\(C_?b-8HbNd04c7XaW]@,UN:RT9C&A]dD^@CCH
7CaVL2(>N3E5-LO.g(I,IN&(,7H(\d2]FadDDg11S8N8gM1Df&62+:=^O]aZTMM8
D?GP(5SV9(]d)G/_SC(#B[4ESdbgONHE,cd_f+UQVDIY]8>ZE-.>SNF9F9EL8FZ=
b(^4c[4,UE:ZW8gB5M0V5,MA=.B5#80\0[95#EP9;W&U2?\d867F7[[9b4d_?cDZ
b42eYJ@+cXRaF=^5c,I_UVV0-RMe)Mf.L>d5aH?YeGTTW2WWX]?E80R.DQB+ZEQ#
F@=^b;1[-1R9D2267]+UAdW2<Y]Y46M=X7eI?&YbY6GeFQ4f.Y<=&=6cXM0CH=8;
fbA5,C,N&\N2WKVO9geC2QX&JRdV<OI^6G[)[gM@^Y/5D),a+2.dDQLF2dd)2FTA
4K:V=><REEP@MS5OUA1,JbYI/XFUMWB925J5XQJQA:QU?C>bVAI74\1aH\e5QM/?
SBFb>,)Y9dI9H?5:XJ;M,CIJB?Hc_V^2WT(71UH.:>3SLNeFUa>(g4G7DHM1@deX
(-:\H<cTb(_O]5DIYAD.4\ZZ\973@S0Ng16E58C&1LeBZUUROR-C?=ES97=ADA5F
IKe9W:1JA7O_^B^KG_KU/H(\8[N+TGYL]/fDG2,fH5G2Va)VEG<OA=QP(A,^BT;S
;H-dfcJVAZe\fEWVQRN]C<]d3D\BCRed\I,MC<.fW=BJL^P=2RC#b#I[=Qb>_?We
[@Dg5\EU1+H3#C;P[c07MO+>20P&-Hc;Z,RP;@RGB@bgD8=D@63.7W)cAK_BW;K7
Y0Gb7-]?_V?W9e:C4V=.6T#@fPIaY=N8()2O)Jb+I6CGY^3#dB<K#/]aB?C?L2c\
+eY?4Ze@.Wf>;eS8B096.0@.DW?\TS97T40-.^AHQ8ZNHVUTIfMRE-PD)?^AaFc^
W(2;8gaS#Q&fWg3-(EUV=ZRJ?+CQ6aJ>4T^430e#D\Z8<(?7UUSOe]_0UEOa(F43
N3E(BWC_5e(d/I25LF:1PMVZQ+Z/#1EP/Q@4)]@c=U3>[:4.[a)C,MRGabCX+ARb
W&VGg:PGX(<f)T#gL<9;-(UUB#)_.IL0G+2S+[&CMV\[(_AfQZL)bDdWSF,-6-He
d3a8cd:2,,B8;dZ##Tg^c56QVN,SB.\2W;R0AZKdGNFO/He0QF>Q]b1cI=KQW>6Y
6CbT(R;-OLG.fM4,T]XcL[DWOCBJGOV_YaR72O81XZ6\#U&eXJ2Sd&?62SWX:?\g
EZJ4BQR9PPgWX??V,XE-AcWS<Q9(/&UA/d1NZ&N7\IO>/<[#R60T6--I,T_?UCE4
EN.IQP/.>-5Ka+RR91Ie1XGR[Q[8O#>8Y[0:ZO?ZB)E=UIWM.^Q44:YCg&30:d[Q
6e)T4/IK;J8PbE9^+<g582W3#MceLeN\cAT_Gf(MSJG^^SgJ1AIO4WQB5X#gZPcR
1F4D-eO;BQQWMH#d5e/C@6eg,/+0@f^Rb<&N.+(K#cIE#\/b9=a8X8O5^[<-+T<?
/ZMAO(c,O0GA[0=1bI))D_>MH-I>M3\.F.?bI)<^+-59(9EAJegb18Zaa^\LUG9d
</V<VROF=NCYaH#HPEV0/DFc1N1aY9[RBSUE0F2<\XJ2YN;/C,Jc-8W:a>U3>0.E
FCXQ\UBJ+CQ]_/&Q;dXKc[KWdAbbW39DQ/2aECC7=1\\fQTTLIf8:c_J)?D^fQR/
cP5@&(6AP6JgeJ8]eN\WXaJ(455^#2](2<F)-70K+1UX<UYP6ILYNZ<\UMS?Z80g
L0S.4VcHcR6gN(JSc,I6)b\A5V+YVeHD?cDAG=)fH6J_A@gBNY&8141N._5]_<0.
+<ES@8F;J?=^fFgM.2CQ2++5_]O6SP32;([QB/-G7e7JYL@GBX6/dX>W12HBNNVG
?FBKK&.ZSe(37_9QN./d<]/[MWfUR#V07:=U2E;^?0/[g-[:cJ?b\Q>cc6[+5J0?
bH)UN;V8D:F#fe?VQdVcN<4I55eC1TK@M1/9,WIV8T53R1>,5gT@CZ6Gc8MN81cV
K;//J]6)#b@aG,D-J:,8aW.^^cb\UCRK71012J?XICA:1#T<>4@6Ce[c#MKC@]\_
86LB,TT73R^g8;JMDFQ]:Cc4:Ca7Cb@>/6JE)PI2H:BB;<\:_8_-/fg)+fGYV=^P
^:P=NN[UdFP:_3VKe.>W7Z24,OE.X=U()HHUd6PW]++VV.a:D4AZH6.85_NJV;/=
UX&+&H@aO(UQMN_S@fN7?AT>fVY,cW;I-a?4<Da]e]ZUDM(#O/6OS29T&@Cd#GC1
?)RL-+ZaS/^/fW+/_T=GL//AMX(BDdfVfT(D>Yf9R[_B=/]EfW(,^^#47;W_bQ1=
,R#L(@XEC(;#_PcG?3\DD.)W;CLY=HD8BVPLLN.[3gQIUF1TNK(_/SB.PG6SZSAc
df@.Y64M:FE;YR0OM[fL1_7.M2GG&JXXYN[GC6,;/)@.99/PUD5],EQXNYc(9;&^
J(/45eL0_F>PM\QM:JP#Xf4M-Ue<Ve6+-Q1T<(.f47@VJ<5dbE17H)b;1VK9a@Z-
]e5+f\OIH/SNA7V<X)H+Z8I.:93UY8FI=CFH>)G?KG72MX5H^EKP?dF/1U3Yb5?8
BE..>\G]WIJ?F1WV.K[aN^b.Ze3RO;>,;b5aPZAJN3>>QX6Ne#.cW9:8b]7]+c=3
,T.ea90KKY(1D6OfW(M/I0=,V[(4SZg[ZA:.3P7NCFDS-1-eCMA\>FVNU&]dBQY;
gJ]-+.c)d@4\cE56X&dXbCR8_ANbLG0.0cCQMZ=:<?KKRL5(LF5Y.3,N:d:c2)[A
V=7AY.YWZ2I19=V1Dd@82M]fC_I9VT::PV02@K2(Ocd:::CL:SbSIKc.KYRE2JM/
9V]bAc4fM_;.18P?HZL&LVQ(PY3YH4a@E<f0JCJ2UIL>gDEE;,gI0UU@44ZHU3[P
V_@XT<5=3gW5d=B@bfN3?@9<RQ1<\g1LAG5bb/[VZa80TLQb.+6^HEc;D58+P-F-
1SI8.fG?SOUg3dPP0?WeG;8>6-1\eYGQA^50Z\5H-7d.XN&^_^DQ3\G<+WC7R5JL
AE.F4E=.P],W9=&D);EM:TLL?[\H?A^_D(5VHIY0[S<KeNSD:K[8YCZ+G\E&LC[A
afg&=YFVR7TIJOO/->O-<(D1Z[\A]gMQ_1S2/.ZOR-M),PL25#TTb=K-JV]7gdKT
<+M7?e4CU:9SPEMA+Kf_,BAM<H+dXP>RDE#9g.g6E_\\0DF[I)/493,,f,VB+>c?
QJ<3-E)+M\>LTc^A:D3[HO64;Ad2YA4c;A<aO>62d2Eb?I_>^,GBg;_VWQDMI0[K
D8?@9gNZaJDW?bF1&4-(R10gaJ\0cXFDI3bO-][IX-Q-FbSV26dI/H=5aX?U^^)R
,=0f94FGQUa-YG>J5#6[</3YA[,,C,(?S)W[BFH]Y[>W;;-A0C@>BQ,PM7(Y@2d/
?Fd8B,VO9Ldd8BVSX#JF\C9P&X6B[Zg=eK)W\[D9M8?eDDRP+K_&()(1YSfTC:,9
+2Xfc488+bZ8c4XSZ[A;E.OG1<4J_+XAg(dCMN#2G.f_6bb-TPN<c5R[<Z#>.(f&
PH<S-HTHJ9\5V+V#/>6LPE5@@NR5T[OSgSRLJg_/?R@_A$
`endprotected
