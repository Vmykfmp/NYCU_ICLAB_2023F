//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Tzu-Yun Huang
//	 Editor		: Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_DRAM.v
//   Module Name : pseudo_DRAM
//   Release version : v3.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_DRAM(
	clk, rst_n,
	AR_VALID, AR_ADDR, R_READY, AW_VALID, AW_ADDR, W_VALID, W_DATA, B_READY,
	AR_READY, R_VALID, R_RESP, R_DATA, AW_READY, W_READY, B_VALID, B_RESP
);

input clk, rst_n;

`protected
d0V12^V\9?BOQ9RN@RDHED3B5TI?CDg(DOL[V-E:3>XBdCNW+2B/.)FSM<//R\K:
0GfWS3cKZ:+9,)eb,A[)UfT^(7V9a;-&eKD&EYdTO?/BB$
`endprotected
input [31:0] AW_ADDR;
input AW_VALID;
output reg AW_READY;

`protected
V_P?dEI-&U[>;?=Z[PRIC3A2<6I>;69ZXaMbWgAD9:I\K)_2Eb43-)/#XeWJFF#b
Jb5NT)>QZYQTT?#&]6(Yaf#X#2-d>IL7?$
`endprotected
input W_VALID;
input [63:0] W_DATA;
output reg W_READY;

`protected
-QJ6A5L,g0@8fQ4R8.F9_WJC]&@36NK9MFH(Pgf#8bfB/7=6,MN&+)fS2d+1G4YS
J1M9G38R;ET.BZN#aLB4Z0@,<7=VeJ=I.BSH@JC;D8IBC$
`endprotected
output reg B_VALID;
output reg [1:0] B_RESP;
input B_READY;

`protected
1EeM\aB,N=B-C)_+@aXRe^.621/I3PAGO:<J+DH<-/T-)I\D;O0F,)b7N^Zg\GQ-
WRe(3Q<(H.@YE/HCQMY8FR4b/1GM[&EbT+JH@FWCYC--A$
`endprotected
input [31:0] AR_ADDR;
input AR_VALID;
output reg AR_READY;

`protected
aC4deLgLWNI#L7-@eJ2E:S;<[4&5WL[.0[Q#XZ1I?^J(E?-;Y+c-2)d?Q]FJ3;1\
VZfCeIM\)\[4:&@7f+@R-)4_:E\;Gd:A>$
`endprotected
output reg [63:0] R_DATA;
output reg R_VALID;
output reg [1:0] R_RESP;
input R_READY;


`protected
-GNB+GcFHQG;ZWFB39<5KI>6a1cc.DA^)[7=Q<HE51W0EX;#WRJc/)H[49W/ZF8D
+][[#CZd@H453EOI,@7d:D#ON7D11<7B9c+\bfTgU+,-VPNPe3(BM-#:E8U-V,bD
5NTTa?RgJI]>Y2=;?#a3W=aP5(\g1PF65.7Lg0G5::A;f>-B42YGL7I,KAS.B587
I:_6);eI1V@S1I#dg_4VM+]Z-1Uda,9&-XOTgGUFR0YO^P6T::8Oad1eZ(N53(8E
EJBV?3f?M#fVK2aSS@KGg\:ACNV3?<e#P;+(R6#QJDE:6S-<Sag=dD825?&ES&g]
0?:OVe;]gb/c&#39CZc_+X/]17+5<AH:c,:\1V]>5bSOdT^9F;9OP?43WA=8A\aU
^[ST7?\6]d#VHAgB:M1KSLPW0ZY]fSH1T_RJ>-&.<8bN>8+32)PWBb+1X\B7FP5B
;aW6\+f18S@NZ>)5SGH2MA1&g:TB/a1I86HX6PdUA]9df+VdLEKa7Yc8LX8EHZ>V
^]XTcC+N&K>@Q]8K85]+NQHTF3Gdf5a>KM;XMDTL8cQ2dF7gV\GN,>Yb8JeAS?PU
F);aOQI[V3,eEAd_afU/bfK^\0Lb.C5;1;]]bE3\(TN(Z_.B<0Qa5gGY3_+Q#1RQ
1/b=EMZTRd]OG[e,NHd]9UB_QfRQ_L38Ba\3D9LQ52EI3Mg<S<0:Ugf^BPVf9fTV
c/6I+PXSeCI6_OKR+TP0aL[O0SRIF;gJ--I^;5V(HH.99ZE3eN@\J]aKFR1LD<56
^1LIc[3]IJLG)2[bgQREdEbO0YKFR<8D.]HV=:U04P\SA[LEX,Db_V4PEODe#CR#
b/>@1WBA,+dSePZ;=PW0C-[9:]RF^&RB[NAg<<F0;7+T/-?A>J&)J>B?.UbL3=?W
9^d\L514R1D<]<FN0)eN?X-#_[:>0geRE&R](Q46C+_OU(SH)Ma2]SEXg(N=8/0X
-f>58N4A+J14f\7d7e)6OTI(C[:TD(?3,,Me53Sa5@-;M0E+ZH7WHAJXV_OKb5:Y
I=6YD3=\b=XAdf-B,G3&M^&-C74[VY7ca]&_IV]5&CRR.2C([1;[&D02)^3Sc</&
Ne&dXJ3R(g:+DdXI0Ya#T30BZL2>2SfgOM5ed[Q;(._Z4R4c&A#HeHDL^\#D9Ne<
I\03J@0aR,[WBR(BY;RL<LKF@69@=F_KZcF75bPZP=V)/WP-_JXXI^g28BH_-BEZ
W=6bVLA38P)12DX<UNK]53^YcW/4]#XZQ6(;]V_:ELK]]I[WcR1?)fbL@I,J#11(
I[?Bf_5#R?R5&NM_Z0G2Q67#^JI=f=ZL1KAMB&HVTY9S>[9O\&d&J00JC5JO8a>1
E9,\J8TYOSL?J<[3(^Z/<(MN\(GFF6XNV8Lg&39U^#H]Td#5D08PG4&;LA?&IdG<
LJZ_ba9+>.XAR([N@gBQ_,CL>I,#7-;&?ceL:a)E\A#5=6CIJ<Q?c-6Rc5KU:DFI
<.U+M:/eJWAW_UVH:9.FKIc,,M8J^;:RVMeBS[8R+([VB6_1PRcH@HP+2;>6g;;R
SQ74)KR<6)(D@P_)DPbPN<fI&S6IXD:@;-2aNXS_W(FaWLW8c;RVec-O0XC5O,=7
W2.Z6[d;HX;B@B_dMDSI;^;<,0cNBFb4geRM<\EYF6M6,cgORg&LbL;R,?3[Q5f/
[@;R^0[Z=SZ>Fg37NPO>2A^[KeJLf55d?+,1.PGE<(3gP./[)^X^DTcCD7DFC?F;
K1db\WcG/<UW==N.Z\;.9_=[\Wa_XM=/b@TS&P#BY>P(7QZA<58#NFMED@P.@=EU
KBY]:YbZ01057L#GUN3R#bZ#51[=bL-Fca_D5Z1=E?5?2g?(JYV^2\c?SE6;).>+
b5L\-P8\Gg;)U)BXTI/]^F06.dCf-e-3O^AP7IN_E8\,^QB:.eURLB+1P9I@CE7Y
?N\T]>1Ua-aKL^1:B<PQR(0W0A?J&DSFVOD-[]2aX+].DOZL;OJd\KVb)f+<,[f&
88NdMQ1cCF-5MPLWRgcWD.a(<aLT++#)PCMUF<\6YRZK&NPT&Y+9:g28&>f\I]H&
3JCgLA&2ZE3aYO(]dKcc\8RHQf+-T8DAe\RM59LIU58^LUg=ZW1:QFN<CAL+9DX2
0N<7J@)Ha?U_DLdI33BeE0[&]GObMA&77QUg3AHGf24Gc[ES;Jg/eP?g(Q@;3;NF
M.VcB>2@NKN(Z.bZ9S?K=6Q76JGLWR#AL0O,-:b&29e<0HXA8F8IP]<DQ2Q=NWEE
ZPDX?M+84.9MNI[f;ac+<C>8[KN25_B7_59S\53agOc;.&4:N;=,+EDAC7,fKL>?
cXK>_9LW1c:&@=5POQ:M<2=dW4;LT/>R4f(#1>]S8Q&T2(a;D5<RG&TcPH+&<X<&
;;GP_T=-]/16[TJW\[;X_A]Y[FY8\&CaM?f^8@.\&)C.RTPWgEF8OR?GN#GB>)GL
9,H/Z<32A/Q.1bYH5Ff_\b4[-XE<H]EZ#Y@JT?820E@bB<Jf,Qf<?)]YD?F4?(X7
Mc.5ZM-UISCK02[.0#BW7aD&GXDb^@=1B4KTOPJ<Y.A?c2CUMSLQ.Jb\\ST^&.GS
25.UcfCA>CW44.e[H?<F=K9W&VNTUAH43bJ)#B9RM,<>E&;+=L(,#N;KJ6<JUU//
981020H,1G+T@GZdfN\9Qa_aVZPbD&gPRG&LQWZ/(THfX=NQVPI/DY+C_:FgbfKa
8)T9#DcJJe>D_BcCZCA?SW/1/LEc\S>@R\VN+777/F(eNL;K^-bBOS.WI\dJ](1W
#=?-YW-I-ON5D<71EKR(1@:d/).C&TC\8FUC8gU#1D931)7^@,IB4N+Efb:MPG;F
85YDIWMM-J4cS9L:?f=RXPUaZS@bLc@(&1N;gCaY-7g;XNN?R5ION#CO6-Be^94S
[c.fI#GKIRSN]D4R<HZ<bP=86Ja_&<.f?-?]>&1cSS)M4]O9dP^5b7>fZUV^YgL\
fEYK;c23=88K6=I_CR+dN-cSf]=-M7I3AJJW:))X#[Ng:QB[LB#CB+AV1g+S1ab(
B>UZYJN@(P+2@C&eH0KEC.FT0G;)6=dJeZ?<,W7C=L[N=]+LAAa&168=#)O_.W.<
-B,NeH[UZc3CTZY8\F8.0fXC[Q48LVKRC8T<a-(D_>/=Tc;1#197CaRZRF)CEGMg
V<0)2.b11I.W#b<LD9UWdZM>M[MB3cPH)B;bLaI^FH+2g5;CgPF^F1V5e5PSV+:H
CH9R=H03N(9db3<6H(:JD[Oc?DbM=[V:TZ#d8C(:>]O3])IDB_VQJO#TC+Z2J</M
=@4BN3_HX5M0c@aTD^PH?(>cM(b[]V4T#NO7QP?;d\TW;2^3(\1=PI?GMP\=6.=?
.H\eE9fB6gG7b0aZ3LQgBO,3X8B&U]2>YY?MM9MVZSP3X=Y[#UB7C3/F2-.9@21P
R:WQ\cYAf-?g]=:3LC+7-WZF9/,SP&VQ3)?fOY-?I=WVMc(VWTL:f:O.VK7DB.G=
[e:0=&NYGPDg7X96)#-(@a<M2E\dLdcHX7X;D6DKKabT@9I2@IUCf/0bOEf>aBJ1
CW:TX=UJ_2=]F&\bfSR_g0H3/2)97S^^^Df=P3Z4U[aWce8KW.T_5#EDIXDOZ+Pg
C^>[3S^d/=FG(C2C\([W<C3ccaRP.d\U1S]=?W:J3ELg_#E9R&K-ZHLa4J;\&a85
0-e<E\(:P[^Oe-B/ZY3bW>40HYQ\035QC-[)gKZ8070Oc<B(D^&WCX4)SA(85[2>
NMO3,FY&IB]\CadS6LIH1985b9Y>T_SLe#W7J5P:aaL=f6#I#;I<_cT+&5N\f.CQ
&MWCE:2K67L__PCBA-?T6XN-g<Q.E/\YS1GXF&[2a_>KVGCKXDRQ]W&e&9KfJe&U
M=U8[=[D6DEg;f^1X]=_^_4Vd(Z1]08?M+#S(Q]7J8:E<^Z):.).YM=L[LN-f5AD
8a0+c]adSL:BV^?M<0bG0O?1a^15>-4NSGP^MM?0?F^[#dQX=K(HZE<KP,JBR_5X
KZE#4(ASDWH+Q9>,8V7TU/dCY^D5-N[^0B\?>RM.Z75\&T2f4_>.W0+.C:L&])IK
KdScB]N>cgM3;Sc-A&4)W^&5.#Ed+91QXBP]2(@U6V[T5Y)+457C,QbT]QW;<:Kf
?<^7/A+.0Pd.N6=QAb>-9QEY+019510e-+]LK33PJCNRKV4XGYRR:A1<&CP)YJMc
dTD9+fE<a)8:ZXHW#SP#NUGF;X&8UKQ,=^RJaf3NY0THXLCUCSaF=85c4G+\3H^R
PR.TKB0X4JH:/2?^ec1=X3C<^HBO<1M/I1?<CDUU=JPf#M9dG@XVXe0#^D@4M=#e
09YTN-fb8)H2c33[?+9Y9bYCC+U(-1c^6E#2e0U+BfPbL/3c\a8H3_8V+)BW0Z6#
(eL1,FH.e<LL(<\WGO3aFW5IR,P>Y:8.K:BWHW)Y#>F=+]>K/NI;(I@<\M+AUM49
Ag,W1=e[dDTLHGcR?)cKcH9O61Y[7gF=^?4Gg8eI__^1^E(0SHPL<CAW)YC7:fWP
6W8_LT/DZA=M_@2\FW<7cUZS3\HFfU4NNI&SG2L4cJ>E4gaPQ;GQ?TbQ@SR+X\V3
=)P6Fa?PfR;EI76K\cZDT^DW)\]eAdVOK0NI1HR8[3_fG:J1Ue9DPK4+\GO-E18W
==RPABc1KI7P#Ne^2c>AN]_4;\H(H)eQA:<UYOWc2^/22-D@O)YT=e;OP>8EdSAS
b5aZNGTZY?3N]J3f>4#gc\+bb6_YQ;[1QR;8[a4;+7UAAR;&8WADB9J7YE#?FcaV
ND<8,1H4EfO=+II\ZIJad7PJ9Z]V6_./9I@S]ad?cJT8]\c9dg/><0\JQWe&83=\
@Z<gaEOD@ZaGE51K\C(B-RNRR#D(/fRH@Y]Y;985d:P:((+M8f)C+04BSfL79BeX
1Tc.BQb6b+dM1OUB=O+TFO12Ne0AKY#S_LCUKC@C6d6#4:B8G,K<B@YFJRH#WP85
M.5^e86A1CGa=Fd1Q7N6V/.U[#?S)P[&3Ccd]/@8NH<=F&<0&;ZLJgYFZFF:YK6f
32&;7T3<UH_#a#8+(XPad_KA.fDI0U?M(XP2#30]T8\0=f=SOMANY@:M9]8J/)OE
-TW(\fLAVY.[\eU[>A(K;0e(^IQ@I@;dK?M]2f>5^Uc9]:+96VZ6P+PO(aE6H.05
KS8TP<C)g]RO@9IF;C+SJ=H9/688(/MU6a2NR?5EO)GdKaV:cJ;Zb0017J&_?+Ve
0]5QL4?C348(Q[^JI>JE[Y9PCQ3c528DUGU[>a)>@?&gfOG(ggM@>a(8deK:K5cX
6?TME2?MVH42C[,<V2cQEW&CK#cBCXH<DOg[]&Z\=fU\&6IQ_U4d7;BL:T/8E/]?
cEV41YG8dI)Ng=V.9f6/.M<;2#BU\J<7&/)=Z-;Z0J?Kb/0,B[K+.ZB@._-b7Nbf
9<\H)[IKHafT:68(Mb&VL)WRN;A&U9E]\B_Z=1c@]Hf/6K7VN>,WBXDR^1;6<U@O
bb\b_e=(PVH5LQ=dMY2(5P9fV;E<_Z)NFO^+[V73.E00PeeHHNLaHP]1J@4J5D&c
e\Q#BfT]8Q/4b3KM77(LINK92.S6XIF\D;7?ffXWVY^1N39AHWW7&2X1T[MS<J6:
fU:4-SBR.<53]Gg8OA\-G\;[UW@]ZC&c:@-&6ID;.5EBdLgFc6YgS^.1P8PTH<IY
ARa^8e5X.-7-;GeeZJ:Teddd.7;IDKF0AOL>(718MK#XD3,B0V5:dBYS^H_V&6(D
1&V&Y/a(^D=g/S\L/cJUFS&Z2/HO@67;A<)FbPTa<faRAb4S+KdE,a,eC^K95@[4
Td8dY03ME=_I\_I<MPF=ad&,\Ca0:(d4c1W3\Y?./\FPV(1?,8(IY/5&()OaZ\..
=6\4H2d6R=O>Aa&YI??>BJHKdE<6PUP\S0fXc_e=I?,eUg14a5b#XT6]8a(QfJ(6
HZV#cABE(C8_6;3+DQZS6AAKK0KLS,eb:c5L.g?DfFZG)+B1LM;5];8:24C;A5I(
JG2P:I4;LU<U]Fb<ZOW.6</D=-Q./52VR4O[\8JLSfKW.O.?Pa<4Xb=T-N)Z>.DE
Y+^@0#\Y7?IeAJSAe]?IH@SEZ8LWOeH98cYU9/fH5FQ0STLY91:ZD;SePBB/[4]H
9WV9fePcFdK(M;T1[ZCF4#74RcP7.&X)&E>171;U9X<(<B@VY\]2QELcRAg)gG.]
0<b(fC+Zdc.:/)Od6Ca1W&:4d[eD49dTP[Yf&f+-,MdHHM,H6BBfF.:89c)0Hc]:
755\JaHfb(B0O?[@5DV7VU[g.\UP_HZ/a?d\Q=@(;-0Z-H_aY3WfBA4O\:ST2G?T
>;9f9B)WW#B,]E+BO4JTPG)VdOcM/9R;,<NWEEA6-IG18^/A-YGE=P@5O[aPTA8g
0Lc9GU.ZGH^C[=K=5H/SZI[\I1G[B]?9a>OaQSOSeWeJMA04LCHd=B&-4HKJ))Ce
3d0cV@ffB<PNM(QIA#P53ON_#ORUe,M[W<3G-\Q?^2Y9,:g]CJ)P_(,/L)1O\.:_
CTa]/_SW4VLD?SX>/[[)aTU+H5\-IVae#BX4R[QN&=e.CP\7FL;8_UW((NFD_DC\
E+NSKIA_V6bAKV?MYR0fP7YWa]L0:6T5^cYafFa^V@^T?XSZ6f@=14Y53MK.D,:-
B_H>Q87+>BbK(G63c@2aF>gI@Y]8WWY>)?7AJZ^_,H_<@M]LgJ?L-SD^U=\/<g>]
<)C+fRB(J.^+C<UH(+c>B.84H.bY/H><46/^X4DEf/G>FT<2eLg+&a.VDf7Cf[^)
HGQb.;X,Q[4:&aa(K@ABGRNK3AEPZgOI->-@U4BP<]>I;baV#P^1UV<VdOX+K/3R
ff13R#+;F_U7b+AE>7He(B7^bPVD[-W[<D.RV.OR^=a]ZX>gUL@/UTUP6?CW78B=
&C22XRU,:^:9gR.[W]R>5aEM>8Z3;L]d^bVHRFcAU0I/NJMWALYaLLRHZ.<1DZ4U
L7_3SdX>eD-G3J#Y-IWKI,DR7>NED4aVI\GV,Y\P2N3gI@A:&\c4,5:aJIQ0\QH[
XIJ?Z_+>-Y++]J=Gf>T/:>b]E7CO#^12PVe)1G#Z.&175acJe--TLOAWB3FU=\)g
Y?5?bQc]BBAWG717_]C/0C]CWA0EMN<G2H/OQ(+?71OS;TI00,1DdR(3<.A[0.#\
+J-9dLJg@)I(14a-EU#4OAMI])[e/2U<PE.J.PI(,1#&;F,L\]69J#>a9)G?<QG5
(5AMK)MD#EMW01=?J)31.VQ0dEMf5#-I78O2E.YGCC^PY(2J5^=68-HU._4Yb9=/
=B[4/f?145W?9dE&#]d/<4Q36;d_b[WSWBGb+,WaGR>LC^Eg8EJ,gV+V2-1M#bI8
.V0;.RJ#C4UQEZB^Z1L_B)gH)b::)1UFY85c(==1D^V>)HVX2CeITG,e8S/);U>&
6#:RG9X]R0X_H>,X=J5BHH-NN-g?-db;B-Y8/cV@^]6K#TWP^4?>A#KbGC^V/<2V
?U?&>@fH)N^6>V+YFbHP&B3_2&a.-+MVZ+YU(,)+>WBg0&EV.-Kf<8_3IV[((Pg&
C8?DP#K<]I1+Q:,LLAUb-#8e+\\4W,-fFT-Hc?RD(ARCSKEF,/A<&QaZF/1Z5>^I
D9:+ZFE,6fb[8fPJS^V9b-X>=Z9&GTgUPZ:46-:Y4EcLG=PV3B0+K+bYFe7WZB3G
WAfF7a-H:#38CIad.#:@(BdY=NM+Ug@_PeGQ5df8^Z.@>;9NQX&La)3MbYSQSO^@
I-LQ/[;N(WbRd]A<Oc\GKb18\<aFK3M7K;^=5=,6Y.S67@>(/8E_7-L@/,<#,O:]
;\eOGPd-MBgX?:IeR4LZ?2QM6N5;@:See,6OLcL7I2FR3)eQ&2OZc]T3-eb&3#EA
L6TMXDUBgcE=CA493V[V9]C4HM)_^8K(C3V3Q6)HC29UR#3H57)8JST2Vf=1-C25
;(COXB^A+Ob^a+IUR_fGHU=ZcC\S_LPU(RRF-Z/)a4d<ag5b8(39L6^.0B=g0Rd8
E7XC@_g&&<:L<W,)?:^U2f7)_+#?,JFKI3?QJ1QV#;aDLW/dKBY#5b)7V/:V53J9
3L@a^,#/2T=35Y+Y><GF^R,T@LG/aJ98=@8ES84Q8Ucf#G7:D9ORb(gBJ#C96gaX
Te918\Y+U_>6E,eFXgTI2))dW4PdX)F9D5EfJVT>TP_;,SR_07afbB7B]#U9T5E,
@3HbSD3IL1B<#1;DD2^fPYR<SgS=BT9WZe\,eSNC=a[58dKV@^/Z)>[/C1A(EU,(
]2_G8W\]FD4.YV<<D.2J^4OK]b@c.3@&1<\-:@5]bKRG0&Wd>U&X1JN&U+6069G[
NOdT;70TE]9Yd6T1-HU,XC1TPX??FELO<1YH,TLg6?L]91S>EC\/XD_f:d>UD>dR
2UCZ)N?\-A;;I4+2e1c=)/69B<8+A5U]-&O,CcNJOP\UEE2#\AXAQMEW3DC61Pe)
(6IN\]03@g])fL@ZHc,bELcV?M,;6a=H//NU^.PO=0Z8/UUFLH=aU#]&CR=fD5IV
+c[8.Rf+#WW>9^40#P9VJM0F+5)AQK,#YeYe:>R7#G.T8D/dFbL@Ue/\Cf5]PL1<
D8ebY.X_5-F=,@2Jf?I8fbPP.^-9NBL=2CVeV\NG)ac@78M=4_AgP[LFAQ/[5GT6
.@8eb:6)H9B3N:3SVg_-]HUge0=7KCGRCZ@M?0ET5-Hc_a5MNe?.Zf#QT7=>HV8@
&[=W6eW[^R>7/VU,RYf+?BK=E:H&c>.gPG2;<M<O0IC0)Xa:DgJ1F(HS0MDFMg=b
a>\A<6\];@6DOf(&&26J^[85/MdR)^/XYTKD6f9<G^^)+,]F?-X[0G]I3A\CIW=Y
1?XPUO5^e+I+GE=)1A#YJW7M/47a-U\We.g45X4UH+S23S+AYI7YdFUGQa+1I@5/
UE^/ADe@f+97D3g@f>AR.(L0Q#\P7a34-Q]1A)UJ.W@GEO4_8eO6MJLK#RE-^HNZ
23CRWeME0JcZ,:]T&)XPE:@D6e:=bDKJ68\=OKEZMQ,EZB-50bS(_2eEUKZI\WE_
VC_.7&f,aE4&,]?I_4Yc27HI4C@2EI?aNW/9CHRBY0OZQaYVd]6MJI:Q;/:(KV2,
Z5f0U5FQg6ZH+7+8f7^1N;1Oa3]gTZg,Rg&b]VEQQB=L(eUOHM6JbN;(=.&4EV-;
J.2cd=EPFOeV:(741@CH/X/7AbF7VSb308\88O2]+;>DVEXL<BcLKNZ9Sf[J/OI&
_Y:OFN/C:=:cL.530I;P5<F3&aK8/_.P-Oa-&XXP8XeKC<a;D^HggZQ93Ge,ZIVX
W7RA-UQZM9OcGb>B9[;Caa_AV:Y0ZJURa_/+QBJ\R2e8PM86YKMScM4Q4dUW;GEL
.3UFdGDcec17cG,28-^;9M,1G>Yec+UQ.P7B#7Q@+c;7c_bG<?&83OeZLdL?[FM>
)a&:aG0gVPWB_5)7;Vb/^?+SQ0X4-GbN-UVD.Q<.RFIX,e.488B:+Ff#7E8]FaLY
>S<?2)M64O719,WK7>.JbbFL/YHI#eg]IaDUM,)gc6Fc++2VY^/(7TYA2F^_W[6]
>I3ORVD&:#YTc:&+.:M_UAGHKKT9<AP4b)@1[[bG02>N<@e0XGS\A=9\c+J2WQ.-
AF_Yg32CVYGIb+ZY)b6U8BbLCL?7?XDIENK/NW9B>KL=/KT81+&c5:0-NQ(e:N^1
9I65?I0?)bB9c912c#HO2T)WeS:XF5/ZGC<A+FDX=WBLd?[1[-R(]_0VB_f2Z@Ne
#K]46@NeCJFQc150B&b02-D7=5P=MfB:I0L3NgT4\.F+J([_eJGV;6Q2>OgPO+SP
C@P9g-+Z;Pe->BQJ/\WEOZ?KGTcZGCMLY:I=K3aAP;OZYec,>&3K;fO3YV/,2XdK
?E5ZR_M6&2Hb^I<US>L[>F(EY>eU=LKU@Y+.>H<YUP[:@=??OF+NUKK9cQ,<^0CS
9;0ONCX>QY]?9KD6#\QZ]PF9=T4H^(0DEc:OaLS,/,]PH_=_<7dXM(.LLc,>0SYH
;08L#3(T)&NNaMU-gN:W.9D^4Z)EV3E9Z#6J[Y-;+>?,Wb?S1W#?(Sd40S644?3X
CC-?U2Y+;&8A;3HD@A.C&^X0fO9?X0c7geE;7gNI:U#0=b+,H,cEP4&G?L;,4b.F
T<-V=V56_]a/=b8=a2E&&G[D+@YDY]Fd]/g0;/W=ZU&)^@GQRTV0>/>+WBNC@,SJ
3]Og<,^]RPNF3[B/-5(Y9AOWO\MZ[>b4U3^EW]XaAUNK_=K)_>f+EWT9^4J3<@gP
VCfe\M57DVSPS<gG)QWF\E\U+[?fXLJ1>XMd2afQe]3T5H83cI?/ec\C>YM;<2VG
I_(EZW+YU4c,e4D;CRSaXP1ANDLMZYR(?0Zb3\ZG<6423&;8PcW\M\g9[WQ?cDdJ
0DfI4+:4R6[b;V,g])<W6Ugf+@BCBAM?g?7ZD?I^<KJ/V2,FaY6FeOLaBS77BAfP
Y3TeM0621G:;<^YMBdY,3G.PWZ7GS@1+a2_+MZY0QKKBAM^GJQ9_?QRAQ7b)40MQ
E;=+F882ML=c]b=UQ@Z=g[LH<46,GXN),K2,f/^K<VFC+B4@7/7Nf(,JF1J.a<KJ
fQ69FST?IbY\a9#10W7+3J-?3A&/EZOB;60=bK9>>3E#?W9?C:/F?#_fSBNTFY0U
<QKQ,7gARf[V\?^.bQ;])PA>0aXV@@L.3OZOJ9.@NL3W^<,JEWDgU[SeQ/eXAFb1
ARXR1DA833NMH1;+W@#,4cHF&^:DQLF,gT2<[3R8#]:b:6^X2M+G412,3H5(2Q.C
Ya83HKY(B<)<[+UM,4TaFIHReK2J4?;)P\0GFGdIY9N[@?O>2b#>0[GA_YW)BZ04
2.@25-S3+D]<41O>-0W>J,_BAS/?Q\&793f=-9##e1@LX0.&g2W(OGc/)7Z//5dO
6a_D(L3#8RJ4)aP]+gfbDC_[1:QP]>CP;f>g,g=)2ZO;fPM83/@8EC+gg7f_D<)J
[IXJDDc[(1Z=__DL:M,fg3BSL]f4;S-/c@<(+D+_0MAXJDg6:/SM@NUdScdO&URR
bG&WZMJ6RcEXLc8cX#<=5WAL0_?XI.U\YJRc6]I9HCK?Bd,<C/GW&cd)fEga>\RV
LdM3TDMM-e;f.=.^Wa92H+MZcESFU]=UP:>8RTE&>>5eLJ7BUZ&^1D2OLT5=K<&>
(^=-?TN^1e.>4)3F]_-T-\#KcQ#S-f6LO(+88HagX+C3<E]P5(\A5G#?03W83-GT
N(8X9(c+4Eg:fO,X;,.Pd2#2\TeB3,>OGPX^KM6S.P&Z@.6UXP:-&0PXDK2A]-ZN
SRB[KMMQVA04e3CFK#+^E<BQ@C?\2NVTZ07]HD:AUH;KbVP\AfUZgT<GfcIU?RYb
:D7IIJF<,^#F:_8,3X@OS3Ub)g+c:09N?$
`endprotected
endmodule
